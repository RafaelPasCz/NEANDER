library ieee;
use ieee.std_logic_1164.all; -- std_logic para detectar erros

entity fft is
    port(
        t      : in std_logic;
        clk    : in std_logic;
        pr, cl : in std_logic;
        q, nq  : out std_logic
    );
end entity;

architecture latch of fft is
    component ffjk is
        port(
            j, k   : in std_logic;
            clk    : in std_logic;
            pr, cl : in std_logic;
            q, nq  : out std_logic
        );
    end component;

    signal sq  : std_logic := '0'; -- opcional -> valor inicial
    signal snq : std_logic := '1';
begin

    u_td : ffjk port map(t, t, clk, pr, cl, q, nq);

end architecture;
